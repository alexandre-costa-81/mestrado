library ieee;
use ieee.std_logic_1164.all;
package example_type is
    type example75f is array(0 to 74) of STD_LOGIC_VECTOR(31 DOWNTO 0);
end package example_type;

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_SIGNED.all;
use IEEE.math_real.all;
use ieee.numeric_std.all;
use work.example_type.all;
--------------------------------------

entity test_receive is

port(
	CLOCK_50: in std_logic;
	UART_TXD: OUT STD_LOGIC;
	UART_RXD: IN STD_LOGIC;
	KEY: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	LEDR: OUT STD_LOGIC_VECTOR(17 DOWNTO 0);
	LEDG: OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
	DATA_OUT : OUT example75f;
	receive_state: OUT integer;
	reset:   in std_logic
);
end test_receive;

architecture KNN_arch of test_receive is
signal x: example75f;
signal starting: std_logic := '1';
SIGNAL TX_DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL TX_START: STD_LOGIC := '0';
SIGNAL TX_BUSY: STD_LOGIC;
SIGNAL RX_DATA: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL RX_BUSY: STD_LOGIC;
SIGNAL WORD_INDEX: INTEGER RANGE 0 TO 3:=0;
SIGNAL DATA0: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DATA1: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DATA2: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL DATA3: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL COLUMN: INTEGER RANGE 0 TO 74:=0;
SIGNAL receiving: integer range 0 to 3 := 0;

COMPONENT TX
PORT(
CLK: IN STD_LOGIC;
START: IN STD_LOGIC;
BUSY: OUT STD_LOGIC;
DATA: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
TX_LINE: OUT STD_LOGIC
);
END COMPONENT TX;

COMPONENT RX
PORT(
CLK: IN STD_LOGIC;
RX_LINE: IN STD_LOGIC;
DATA: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
BUSY: OUT STD_LOGIC
);
END COMPONENT RX;

BEGIN
	C1: TX PORT MAP(CLOCK_50, TX_START, TX_BUSY, TX_DATA, UART_TXD);
	C2: RX PORT MAP(CLOCK_50, UART_RXD, RX_DATA, RX_BUSY);  
	PROCESS(CLOCK_50)
	variable y: std_logic;
	variable etapa: integer range 0 to 10:=0;
	variable countc: integer range 0 to 77:=0;
	variable countr: integer range 0 to 77:=0;
	variable count_wait: integer range 0 to 5000002:=0;
	BEGIN	
		if (reset = '1') then
			receiving <= 0;		
		ELSIF(CLOCK_50'EVENT AND CLOCK_50='1') THEN
			IF(receiving=0 AND TX_BUSY='0') THEN
				TX_DATA <= "11111111";
				TX_START <= '1';
				receiving <= 1;
			ELSE
				TX_START <= '0';
			END IF;
			IF(receiving = 1 AND RX_BUSY='0') THEN
				IF(WORD_INDEX=0) THEN
					DATA0 <= RX_DATA;
					WORD_INDEX <= WORD_INDEX+1;
				ELSIF(WORD_INDEX=1) THEN
					DATA1 <= RX_DATA;
					WORD_INDEX <= WORD_INDEX+1;
				ELSIF(WORD_INDEX=2) THEN
					DATA2 <= RX_DATA;
					WORD_INDEX <= WORD_INDEX+1;
				ELSIF(WORD_INDEX=3) THEN
					DATA3 <= RX_DATA;
					x(COLUMN) <= DATA0 & DATA1 & DATA2 & DATA3;
					COLUMN <= COLUMN + 1;
					WORD_INDEX <= 0;
					IF(COLUMN = 75) THEN --75, 0 to 74
						COLUMN <= 0;
						receiving <= 2;
						--DATA_OUT <= x;
					END IF;
				END IF;
			end if;
		END IF;
		--DATA_OUT <= ("10111110011101100001100001001000","10111110000100111110010011101111","00111111100110110111101001001110","10111110011011101101000011110110","00111110010101101101000110011110","00111111101000000011110010011111","10111110011001011011111011100100","00111111000010011001011111100101","00111111101000101101110001011101","10111110010001100001111000001100","00111111001011101010110111000101","00111111101000100101001101100101","10111110101111101000100001111011","00111110110000100111110100000011","01000100100101010100000000000000","10111110110111101011001110111100","00111101110100101000101011100111","00111111100100100010111100000110","10111110110011010011100110111001","10111101110100110111010000110110","00111111100001010110100001110011","10111110110010001101001000011100","10111110000011011111101101010000","00111111100001010001000101001001","10111101010110101100100110110000","00111110101111010011010011011111","00111111101001001010011011001010","10111100101001010010101011000111","00111101110111101001100011011101","00111111101000011101010010010101","00111011100100100001010001101010","10111101101111110101110101111001","00111111100100111011100110001100","10111100101101110000110011011101","10111110000001010011010111001010","00111111100100001010101101100000","10111110100111011100010110110101","10111110000010111001011001101100","00111111100100111110100010111100","10111110110110000000101101000110","10111110111110010011110011001101","00111111100011011101110011000110","10111110111110000010011001100111","10111111011010010111101110100110","00111111100110110010001100100101","10111110111000010100011111010000","10111111011010100101001011001110","00111111100011100010001111100010","10111110001000001000000001110011","10111110000100100110000101111100","00111111100110001011001111100101","10111101011001001001001010111100","10111111000000000010111010101001","00111111100010111101001011001000","00111110100011010110000110010001","10111111010011011001010101010111","00111111100000010001101100011110","00111110100111001101000000110101","10111111010001101001011011010101","00111111011001011000001010101010","10111110011010000100011011101001","00111110111010101110000101101001","00111111101000100111110001011011","10111110101111100010000110111000","10111110001111010100111000001001","00111111100001000010011000000011","10111110101101001010000110101101","10111110000000110010011101100111","01000100100001000010000000000000","10111101000001011010000010111110","10111110001100100011100010010111","00111111100011001110010000010001","00111100010110101010100100101110","10111110000110111010100011000110","00111111100100100000001101110001");
		DATA_OUT <= ("10111111000011100100100100101100",
"10111110000100000111011111001101",
"00111111101111001100111001110000",
"10111111000010101000100100100010",
"00111110010001111001000011111011",
"00111111110000011101100011011000",
"10111111000001011100100100001100",
"00111111000000110001000000000010",
"00111111110001001111011100010010",
"10111111000001110100000111000000",
"00111111001010011011111011000010",
"00111111110000010001111110110100",
"10111111001110010110000010100110",
"00111110110000100111010011100010",
"00111111101111100111111010100110",
"10111111011001011100010101100001",
"00111110101111011011001100011000",
"00111111101101001010001100101111",
"10111111010101011001100110111011",
"00111111000100001100100111111011",
"00111111101010111000101110101100",
"10111111010011110111010001011000",
"00111111001001101000111010010011",
"00111111101011011000110111001110",
"10111110101011000010000100111010",
"00111110101101000100110010111110",
"00111111110001001100110000100101",
"10111110000101010010010001111101",
"00111110101111001010000011100100",
"00111111101110110000010111111011",
"10111110001101111100101000100001",
"00111111000101011010101010000010",
"00111111101100100011100111010110",
"10111110010011000100111101111111",
"00111111001010011110001010111101",
"00111111101100100101001001101001",
"10111111001000010010100111111110",
"10111110000001100111010001001011",
"00111111101101011111100010100001",
"10111111001011011000101011101100",
"10111110111011101100010101101101",
"00111111101001001101001101011011",
"10111111010000001001100010010001",
"10111111010101100010101011000011",
"00111111100110011011110000000010",
"10111111001110010111100100000111",
"10111111010111000110001010010001",
"00111111100010000111011010011111",
"10111110111010000000111010001101",
"10111110000100101111101010010100",
"00111111101110011110100000111110",
"10111110111000101010010000110011",
"10111111000000011101110111110100",
"00111111101110000001101111011010",
"10111110111001110000110110000100",
"10111111011000001010110101011000",
"00111111110000011111111110000010",
"10111110110110110110001010100110",
"10111111011001000101100111101010",
"00111111101100000000011100110101",
"10111111000001110010001100010100",
"00111110110111101100010110110000",
"00111111110001000111101100110101",
"10111111010010111010000001110011",
"00111111001110111101101101011110",
"00111111101011110100110110111110",
"10111111010100110101000110001011",
"00111111001100000011010001011101",
"00111111101010100011100111010110",
"10111110010111101000111100101010",
"00111111001111011110010111100010",
"00111111101100100110010101101011",
"10111110011110010100001110011110",
"00111111001000101001010010001010",
"00111111101100101100111001000110");
		receiving <= 2;
		receive_state <= receiving;
	END PROCESS;
end KNN_arch;